Vin 1   0   AC  12  0   60
R1  1   2   100
R2  3   0   50
R3  3   0   50
C1  2   0   0.01
L1  2   3   0.01
L2  3   0   0.01

.tran 0.0005  0.2



