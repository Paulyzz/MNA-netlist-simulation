Vin 1   0   AC  12  0   60
R1  3   0   100
L1  2   3   1000
C1  3   4   0.01
R2  4   0   100
C2  2   0   0.01
R3  2   1   100
L2  4   0   0.01


.tran 0.0005  0.2