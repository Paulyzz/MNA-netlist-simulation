V1 1 0 AC 12 0 100
R1 2 1 100
C1 2 0 1
L1 3 2 1
L2 2 1 1
R2 3 0 100

.tran 0.0005  0.2